* cell inv1
* pin X
* pin VDD
* pin A
* pin VSS
.SUBCKT inv1 3 2 4 1
* net 1 X
* net 2 VDD
* net 3 A
* net 4 VSS
* device instance $1 r0 *1 3,23.5 PMOS
M$1 2 3 1 2 PMOS L=1U W=6U AS=12P AD=12P PS=16U PD=16U
* device instance $2 r0 *1 3,3.5 NMOS
M$2 4 3 1 4 NMOS L=1U W=2U AS=4P AD=4P PS=8U PD=8U
.ENDS inv1$1

* cell sff1
* pin CK
* pin D
* pin QB
* pin Q
* pin VDD
* pin VSS
.SUBCKT sff1 2 4 11 10 9 18 23
* net 2 CK
* net 4 D
* net 9 S
* net 10 QB
* net 11 Q
* net 18 VDD
* net 23 VSS
* device instance $1 r0 *1 12.5,23.5 PMOS
M$1 18 4 19 18 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $2 r0 *1 14.5,23.5 PMOS
M$2 19 1 5 18 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $3 r0 *1 17.5,23.5 PMOS
M$3 5 3 20 18 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $4 r0 *1 19.5,23.5 PMOS
M$4 20 6 18 18 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $5 r0 *1 22.5,23.5 PMOS
M$5 18 5 6 18 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $6 r0 *1 25.5,23.5 PMOS
M$6 6 9 18 18 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $7 r0 *1 28.5,23.5 PMOS
M$7 18 6 21 18 PMOS L=1U W=6U AS=6P AD=7.5P PS=8U PD=8.5U
* device instance $8 r0 *1 32,23.5 PMOS
M$8 21 3 7 18 PMOS L=1U W=6U AS=7.5P AD=6P PS=8.5U PD=8U
* device instance $9 r0 *1 35,23.5 PMOS
M$9 7 1 22 18 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $10 r0 *1 37,23.5 PMOS
M$10 22 8 18 18 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $11 r0 *1 40,23.5 PMOS
M$11 18 7 8 18 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $12 r0 *1 43,23.5 PMOS
M$12 8 9 18 18 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $13 r0 *1 49.5,23.5 PMOS
M$13 10 8 18 18 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $14 r0 *1 52.5,23.5 PMOS
M$14 18 10 11 18 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $15 r0 *1 3,23.5 PMOS
M$15 1 2 18 18 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $16 r0 *1 6,23.5 PMOS
M$16 18 1 3 18 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $17 r0 *1 49.5,3.5 NMOS
M$17 10 8 23 23 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $18 r0 *1 52.5,3.5 NMOS
M$18 23 10 11 23 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $19 r0 *1 31,3.5 NMOS
M$19 23 6 15 23 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $20 r0 *1 33,3.5 NMOS
M$20 15 1 7 23 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $21 r0 *1 36,3.5 NMOS
M$21 7 3 16 23 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $22 r0 *1 38,3.5 NMOS
M$22 16 8 23 23 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $23 r0 *1 41,3.5 NMOS
M$23 23 7 17 23 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $24 r0 *1 43,3.5 NMOS
M$24 17 9 8 23 NMOS L=1U W=2U AS=1P AD=4P PS=3U PD=8U
* device instance $25 r0 *1 12.5,3.5 NMOS
M$25 23 4 12 23 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $26 r0 *1 14.5,3.5 NMOS
M$26 12 3 5 23 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $27 r0 *1 17.5,3.5 NMOS
M$27 5 1 13 23 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $28 r0 *1 19.5,3.5 NMOS
M$28 13 6 23 23 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $29 r0 *1 22.5,3.5 NMOS
M$29 23 5 14 23 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $30 r0 *1 24.5,3.5 NMOS
M$30 14 9 6 23 NMOS L=1U W=2U AS=1P AD=4P PS=3U PD=8U
* device instance $31 r0 *1 3,3.5 NMOS
M$31 1 2 23 23 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $32 r0 *1 6,3.5 NMOS
M$32 23 1 3 23 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS sff1$1

* cell nr31$1
* pin X
* pin VDD
* pin A
* pin B
* pin C
* pin VSS
.SUBCKT nr31 3 4 5 2 8 1
* net 1 X
* net 2 VDD
* net 3 A
* net 4 B
* net 5 C
* net 8 VSS
* device instance $1 r0 *1 4,23.5 PMOS
M$1 2 3 7 2 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $2 r0 *1 6,23.5 PMOS
M$2 7 4 6 2 PMOS L=1U W=6U AS=3P AD=3P PS=7U PD=7U
* device instance $3 r0 *1 8,23.5 PMOS
M$3 6 5 1 2 PMOS L=1U W=6U AS=3P AD=12P PS=7U PD=16U
* device instance $4 r0 *1 3,3.5 NMOS
M$4 8 3 1 8 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $5 r0 *1 6,3.5 NMOS
M$5 1 4 8 8 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $6 r0 *1 9,3.5 NMOS
M$6 8 5 1 8 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS nr31

* cell na31$1
* pin X
* pin VDD
* pin B
* pin A
* pin C
* pin VSS
.SUBCKT na31 4 3 5 2 8 1
* net 1 X
* net 2 VDD
* net 3 B
* net 4 A
* net 5 C
* net 8 VSS
* device instance $1 r0 *1 3,23.5 PMOS
M$1 2 4 1 2 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 6,23.5 PMOS
M$2 1 3 2 2 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $3 r0 *1 9,23.5 PMOS
M$3 2 5 1 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $4 r0 *1 3,3.5 NMOS
M$4 8 4 7 8 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $5 r0 *1 5,3.5 NMOS
M$5 7 3 6 8 NMOS L=1U W=2U AS=1P AD=1P PS=3U PD=3U
* device instance $6 r0 *1 7,3.5 NMOS
M$6 6 5 1 8 NMOS L=1U W=2U AS=1P AD=4P PS=3U PD=8U
.ENDS na31

* cell inv4$1
* pin A
* pin VDD
* pin X
* pin VSS
.SUBCKT inv4 1 2 4 3
* net 1 A
* net 2 VDD
* net 3 X
* net 4 VSS
* device instance $1 r0 *1 3,23.5 PMOS
M$1 2 1 3 2 PMOS L=1U W=24U AS=30P AD=30P PS=40U PD=40U
* device instance $5 r0 *1 3,3.5 NMOS
M$5 4 1 3 4 NMOS L=1U W=8U AS=10P AD=10P PS=20U PD=20U
.ENDS inv4

* cell dff1m2$1
* pin CK
* pin D
* pin QB
* pin Q
* pin VDD
* pin VSS
.SUBCKT dff1m2 2 4 8 7 15 20
* net 2 CK
* net 4 D
* net 7 QB
* net 8 Q
* net 15 VDD
* net 20 VSS
* device instance $1 r0 *1 45.5,23.5 PMOS
M$1 7 6 15 15 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 48.5,23.5 PMOS
M$2 15 7 8 15 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $3 r0 *1 29,23.5 PMOS
M$3 15 11 18 15 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $4 r0 *1 31,23.5 PMOS
M$4 18 3 13 15 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $5 r0 *1 34,23.5 PMOS
M$5 13 1 19 15 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $6 r0 *1 36,23.5 PMOS
M$6 19 6 15 15 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $7 r0 *1 39,23.5 PMOS
M$7 15 13 6 15 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $8 r0 *1 12.5,23.5 PMOS
M$8 15 4 16 15 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $9 r0 *1 14.5,23.5 PMOS
M$9 16 1 5 15 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $10 r0 *1 17.5,23.5 PMOS
M$10 5 3 17 15 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $11 r0 *1 19.5,23.5 PMOS
M$11 17 11 15 15 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $12 r0 *1 22.5,23.5 PMOS
M$12 15 5 11 15 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $13 r0 *1 3,23.5 PMOS
M$13 1 2 15 15 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $14 r0 *1 6,23.5 PMOS
M$14 15 1 3 15 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $15 r0 *1 45.5,3.5 NMOS
M$15 7 6 20 20 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $16 r0 *1 48.5,3.5 NMOS
M$16 20 7 8 20 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $17 r0 *1 29,3.5 NMOS
M$17 20 11 12 20 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $18 r0 *1 31,3.5 NMOS
M$18 12 1 13 20 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $19 r0 *1 34,3.5 NMOS
M$19 13 3 14 20 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $20 r0 *1 36,3.5 NMOS
M$20 14 6 20 20 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $21 r0 *1 39,3.5 NMOS
M$21 20 13 6 20 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $22 r0 *1 3,3.5 NMOS
M$22 1 2 20 20 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $23 r0 *1 6,3.5 NMOS
M$23 20 1 3 20 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $24 r0 *1 12.5,3.5 NMOS
M$24 20 4 9 20 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $25 r0 *1 14.5,3.5 NMOS
M$25 9 3 5 20 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $26 r0 *1 17.5,3.5 NMOS
M$26 5 1 10 20 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $27 r0 *1 19.5,3.5 NMOS
M$27 10 11 20 20 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $28 r0 *1 22.5,3.5 NMOS
M$28 20 5 11 20 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS dff1m2

* cell buf2$1
* pin Y
* pin VDD
* pin A
* pin VSS
.SUBCKT buf2 4 3 5 2
* net 2 Y
* net 3 VDD
* net 4 A
* net 5 VSS
* device instance $1 r0 *1 3,23.5 PMOS
M$1 1 4 3 3 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 6,23.5 PMOS
M$2 3 1 2 3 PMOS L=1U W=12U AS=12P AD=18P PS=16U PD=24U
* device instance $4 r0 *1 3,3.5 NMOS
M$4 1 4 5 5 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $5 r0 *1 6,3.5 NMOS
M$5 5 1 2 5 NMOS L=1U W=4U AS=4P AD=6P PS=8U PD=12U
.ENDS buf2

* cell rff1m2$1
* pin Q
* pin CK
* pin D
* pin QB
* pin VDD
* pin VSS
.SUBCKT rff1m2 3 5 1 10 8 16 23
* net 1 Q
* net 3 CK
* net 5 D
* net 8 R
* net 10 QB
* net 16 VDD
* net 23 VSS
* device instance $1 r0 *1 49.5,23.5 PMOS
M$1 10 9 16 16 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 52.5,23.5 PMOS
M$2 16 10 1 16 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $3 r0 *1 31,23.5 PMOS
M$3 16 7 20 16 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $4 r0 *1 33,23.5 PMOS
M$4 20 4 13 16 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $5 r0 *1 36,23.5 PMOS
M$5 13 2 21 16 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $6 r0 *1 38,23.5 PMOS
M$6 21 9 16 16 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $7 r0 *1 41,23.5 PMOS
M$7 16 13 22 16 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $8 r0 *1 43,23.5 PMOS
M$8 22 8 9 16 PMOS L=1U W=6U AS=3P AD=12P PS=7U PD=16U
* device instance $9 r0 *1 12.5,23.5 PMOS
M$9 16 5 17 16 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $10 r0 *1 14.5,23.5 PMOS
M$10 17 2 6 16 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $11 r0 *1 17.5,23.5 PMOS
M$11 6 4 18 16 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $12 r0 *1 19.5,23.5 PMOS
M$12 18 7 16 16 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $13 r0 *1 22.5,23.5 PMOS
M$13 16 6 19 16 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $14 r0 *1 24.5,23.5 PMOS
M$14 19 8 7 16 PMOS L=1U W=6U AS=3P AD=12P PS=7U PD=16U
* device instance $15 r0 *1 3,23.5 PMOS
M$15 2 3 16 16 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $16 r0 *1 6,23.5 PMOS
M$16 16 2 4 16 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $17 r0 *1 49.5,3.5 NMOS
M$17 10 9 23 23 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $18 r0 *1 52.5,3.5 NMOS
M$18 23 10 1 23 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $19 r0 *1 12.5,3.5 NMOS
M$19 23 5 11 23 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $20 r0 *1 14.5,3.5 NMOS
M$20 11 4 6 23 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $21 r0 *1 17.5,3.5 NMOS
M$21 6 2 12 23 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $22 r0 *1 19.5,3.5 NMOS
M$22 12 7 23 23 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $23 r0 *1 22.5,3.5 NMOS
M$23 23 6 7 23 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $24 r0 *1 25.5,3.5 NMOS
M$24 7 8 23 23 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $25 r0 *1 28.5,3.5 NMOS
M$25 23 7 14 23 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $26 r0 *1 30.5,3.5 NMOS
M$26 14 2 13 23 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $27 r0 *1 33.5,3.5 NMOS
M$27 13 4 15 23 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $28 r0 *1 35.5,3.5 NMOS
M$28 15 9 23 23 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $29 r0 *1 38.5,3.5 NMOS
M$29 23 13 9 23 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $30 r0 *1 41.5,3.5 NMOS
M$30 9 8 23 23 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $31 r0 *1 3,3.5 NMOS
M$31 2 3 23 23 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $32 r0 *1 6,3.5 NMOS
M$32 23 2 4 23 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS rff1m2$1

* cell nr222$1
* pin X
* pin VDD
* pin A0
* pin A1
* pin B1
* pin B0
* pin VSS
.SUBCKT nr222 4 5 7 6 3 10 1
* net 1 X
* net 3 VDD
* net 4 A0
* net 5 A1
* net 6 B1
* net 7 B0
* net 10 VSS
* device instance $1 r0 *1 3,22 PMOS
M$1 2 4 3 3 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 6,22 PMOS
M$2 3 5 2 3 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $3 r0 *1 9,22 PMOS
M$3 2 6 1 3 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $4 r0 *1 12,22 PMOS
M$4 1 7 2 3 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $5 r0 *1 3,3.5 NMOS
M$5 10 4 9 10 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $6 r0 *1 5,3.5 NMOS
M$6 9 5 1 10 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $7 r0 *1 8,3.5 NMOS
M$7 1 6 8 10 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $8 r0 *1 10,3.5 NMOS
M$8 8 7 10 10 NMOS L=1U W=2U AS=1P AD=4P PS=3U PD=8U
.ENDS nr222

* cell na222$1
* pin VDD
* pin X
* pin B0
* pin B1
* pin A1
* pin A0
* pin VSS
.SUBCKT na222 7 6 4 5 1 10 3
* net 1 VDD
* net 3 X
* net 4 B0
* net 5 B1
* net 6 A1
* net 7 A0
* net 10 VSS
* device instance $1 r0 *1 4,23.5 PMOS
M$1 1 7 9 1 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $2 r0 *1 6,23.5 PMOS
M$2 9 6 3 1 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $3 r0 *1 9,23.5 PMOS
M$3 3 5 8 1 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $4 r0 *1 11,23.5 PMOS
M$4 8 4 1 1 PMOS L=1U W=6U AS=3P AD=12P PS=7U PD=16U
* device instance $5 r0 *1 3,5 NMOS
M$5 2 7 10 10 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $6 r0 *1 6,5 NMOS
M$6 10 6 2 10 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $7 r0 *1 9,5 NMOS
M$7 2 5 3 10 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $8 r0 *1 12,5 NMOS
M$8 3 4 2 10 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS na222

* cell inv2$1
* pin A
* pin X
* pin VDD
* pin VSS
.SUBCKT inv2 1 3 4 2
* net 1 A
* net 2 X
* net 3 VDD
* net 4 VSS
* device instance $1 r0 *1 3,23.5 PMOS
M$1 3 1 2 3 PMOS L=1U W=12U AS=18P AD=18P PS=24U PD=24U
* device instance $3 r0 *1 3,3.5 NMOS
M$3 4 1 2 4 NMOS L=1U W=4U AS=6P AD=6P PS=12U PD=12U
.ENDS inv2

* cell dff1
* pin CK
* pin D
* pin QB
* pin Q
* pin VDD
* pin VSS
.SUBCKT dff1 2 4 9 8 15 20
* net 2 CK
* net 4 D
* net 8 QB
* net 9 Q
* net 15 VDD
* net 20 VSS
* device instance $1 r0 *1 45.5,23.5 PMOS
M$1 8 7 15 15 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 48.5,23.5 PMOS
M$2 15 8 9 15 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $3 r0 *1 29,23.5 PMOS
M$3 15 6 18 15 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $4 r0 *1 31,23.5 PMOS
M$4 18 3 13 15 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $5 r0 *1 34,23.5 PMOS
M$5 13 1 19 15 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $6 r0 *1 36,23.5 PMOS
M$6 19 7 15 15 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $7 r0 *1 39,23.5 PMOS
M$7 15 13 7 15 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $8 r0 *1 12.5,23.5 PMOS
M$8 15 4 16 15 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $9 r0 *1 14.5,23.5 PMOS
M$9 16 1 5 15 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $10 r0 *1 17.5,23.5 PMOS
M$10 5 3 17 15 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $11 r0 *1 19.5,23.5 PMOS
M$11 17 6 15 15 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $12 r0 *1 22.5,23.5 PMOS
M$12 15 5 6 15 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $13 r0 *1 3,23.5 PMOS
M$13 1 2 15 15 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $14 r0 *1 6,23.5 PMOS
M$14 15 1 3 15 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $15 r0 *1 45.5,3.5 NMOS
M$15 8 7 20 20 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $16 r0 *1 48.5,3.5 NMOS
M$16 20 8 9 20 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $17 r0 *1 29,3.5 NMOS
M$17 20 6 12 20 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $18 r0 *1 31,3.5 NMOS
M$18 12 1 13 20 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $19 r0 *1 34,3.5 NMOS
M$19 13 3 14 20 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $20 r0 *1 36,3.5 NMOS
M$20 14 7 20 20 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $21 r0 *1 39,3.5 NMOS
M$21 20 13 7 20 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $22 r0 *1 3,3.5 NMOS
M$22 1 2 20 20 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $23 r0 *1 6,3.5 NMOS
M$23 20 1 3 20 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $24 r0 *1 12.5,3.5 NMOS
M$24 20 4 10 20 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $25 r0 *1 14.5,3.5 NMOS
M$25 10 3 5 20 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $26 r0 *1 17.5,3.5 NMOS
M$26 5 1 11 20 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $27 r0 *1 19.5,3.5 NMOS
M$27 11 6 20 20 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $28 r0 *1 22.5,3.5 NMOS
M$28 20 5 6 20 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS dff1

* cell buf1$1
* pin VDD
* pin Y
* pin A
* pin VSS
.SUBCKT buf1 4 1 5 3
* net 1 VDD
* net 3 Y
* net 4 A
* net 5 VSS
* device instance $1 r0 *1 3,23.5 PMOS
M$1 2 4 1 1 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 6,23.5 PMOS
M$2 1 2 3 1 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $3 r0 *1 3,3.5 NMOS
M$3 2 4 5 5 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $4 r0 *1 6,3.5 NMOS
M$4 5 2 3 5 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS buf1

* cell rff1$1
* pin CK
* pin D
* pin QB
* pin Q
* pin VDD
* pin VSS
.SUBCKT rff1 2 4 11 10 7 16 23
* net 2 CK
* net 4 D
* net 7 R
* net 10 QB
* net 11 Q
* net 16 VDD
* net 23 VSS
* device instance $1 r0 *1 49.5,23.5 PMOS
M$1 10 8 16 16 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 52.5,23.5 PMOS
M$2 16 10 11 16 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $3 r0 *1 31,23.5 PMOS
M$3 16 6 20 16 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $4 r0 *1 33,23.5 PMOS
M$4 20 3 9 16 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $5 r0 *1 36,23.5 PMOS
M$5 9 1 21 16 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $6 r0 *1 38,23.5 PMOS
M$6 21 8 16 16 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $7 r0 *1 41,23.5 PMOS
M$7 16 9 22 16 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $8 r0 *1 43,23.5 PMOS
M$8 22 7 8 16 PMOS L=1U W=6U AS=3P AD=12P PS=7U PD=16U
* device instance $9 r0 *1 12.5,23.5 PMOS
M$9 16 4 17 16 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $10 r0 *1 14.5,23.5 PMOS
M$10 17 1 5 16 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $11 r0 *1 17.5,23.5 PMOS
M$11 5 3 18 16 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $12 r0 *1 19.5,23.5 PMOS
M$12 18 6 16 16 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $13 r0 *1 22.5,23.5 PMOS
M$13 16 5 19 16 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $14 r0 *1 24.5,23.5 PMOS
M$14 19 7 6 16 PMOS L=1U W=6U AS=3P AD=12P PS=7U PD=16U
* device instance $15 r0 *1 3,23.5 PMOS
M$15 1 2 16 16 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $16 r0 *1 6,23.5 PMOS
M$16 16 1 3 16 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $17 r0 *1 49.5,3.5 NMOS
M$17 10 8 23 23 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $18 r0 *1 52.5,3.5 NMOS
M$18 23 10 11 23 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $19 r0 *1 12.5,3.5 NMOS
M$19 23 4 12 23 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $20 r0 *1 14.5,3.5 NMOS
M$20 12 3 5 23 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $21 r0 *1 17.5,3.5 NMOS
M$21 5 1 13 23 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $22 r0 *1 19.5,3.5 NMOS
M$22 13 6 23 23 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $23 r0 *1 22.5,3.5 NMOS
M$23 23 5 6 23 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $24 r0 *1 25.5,3.5 NMOS
M$24 6 7 23 23 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $25 r0 *1 28.5,3.5 NMOS
M$25 23 6 14 23 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $26 r0 *1 30.5,3.5 NMOS
M$26 14 1 9 23 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $27 r0 *1 33.5,3.5 NMOS
M$27 9 3 15 23 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $28 r0 *1 35.5,3.5 NMOS
M$28 15 8 23 23 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $29 r0 *1 38.5,3.5 NMOS
M$29 23 9 8 23 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $30 r0 *1 41.5,3.5 NMOS
M$30 8 7 23 23 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $31 r0 *1 3,3.5 NMOS
M$31 1 2 23 23 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $32 r0 *1 6,3.5 NMOS
M$32 23 1 3 23 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS rff1$1

* cell nr212
* pin X
* pin VDD
* pin B0
* pin A0
* pin A1
* pin VSS
.SUBCKT nr212 5 6 4 2 8 1
* net 1 X
* net 2 VDD
* net 4 B0
* net 5 A0
* net 6 A1
* net 8 VSS
* device instance $1 r0 *1 3,23.5 PMOS
M$1 3 5 2 2 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 6,23.5 PMOS
M$2 2 6 3 2 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $3 r0 *1 9,23.5 PMOS
M$3 3 4 1 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $4 r0 *1 3,3.5 NMOS
M$4 8 5 7 8 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $5 r0 *1 5,3.5 NMOS
M$5 7 6 1 8 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $6 r0 *1 8,3.5 NMOS
M$6 1 4 8 8 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS nr212

* cell na212
* pin VDD
* pin X
* pin A0
* pin A1
* pin B0
* pin VSS
.SUBCKT na212 3 4 5 1 8 2
* net 1 VDD
* net 2 X
* net 3 A0
* net 4 A1
* net 5 B0
* net 8 VSS
* device instance $1 r0 *1 4,23.5 PMOS
M$1 1 3 7 1 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $2 r0 *1 6,23.5 PMOS
M$2 7 4 2 1 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $3 r0 *1 9,23.5 PMOS
M$3 2 5 1 1 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $4 r0 *1 3,3.5 NMOS
M$4 6 3 8 8 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $5 r0 *1 6,3.5 NMOS
M$5 8 4 6 8 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $6 r0 *1 9,3.5 NMOS
M$6 6 5 2 8 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS na212

* cell cinv$1
* pin OE
* pin VDD
* pin X
* pin A
* pin VSS
.SUBCKT cinv 5 1 3 8 4
* net 1 OE
* net 3 VDD
* net 4 X
* net 5 A
* net 8 VSS
* device instance $1 r0 *1 3,23.5 PMOS
M$1 2 1 3 3 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 6,23.5 PMOS
M$2 3 2 6 3 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $3 r0 *1 8,23.5 PMOS
M$3 6 5 4 3 PMOS L=1U W=6U AS=3P AD=12P PS=7U PD=16U
* device instance $4 r0 *1 3,3.5 NMOS
M$4 2 1 8 8 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $5 r0 *1 6,3.5 NMOS
M$5 8 1 7 8 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $6 r0 *1 8,3.5 NMOS
M$6 7 5 4 8 NMOS L=1U W=2U AS=1P AD=4P PS=3U PD=8U
.ENDS cinv

* cell an41$1
* pin D
* pin Y
* pin VDD
* pin C
* pin B
* pin A
* pin VSS
.SUBCKT an41 7 6 5 1 4 11 3
* net 1 D
* net 3 Y
* net 4 VDD
* net 5 C
* net 6 B
* net 7 A
* net 11 VSS
* device instance $1 r0 *1 3,23.5 PMOS
M$1 4 7 2 4 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 6,23.5 PMOS
M$2 2 6 4 4 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $3 r0 *1 9,23.5 PMOS
M$3 4 5 2 4 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $4 r0 *1 12,23.5 PMOS
M$4 2 1 4 4 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $5 r0 *1 15,23.5 PMOS
M$5 4 2 3 4 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $6 r0 *1 3,3.5 NMOS
M$6 2 7 9 11 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $7 r0 *1 5,3.5 NMOS
M$7 9 6 8 11 NMOS L=1U W=2U AS=1P AD=1P PS=3U PD=3U
* device instance $8 r0 *1 7,3.5 NMOS
M$8 8 5 10 11 NMOS L=1U W=2U AS=1P AD=1P PS=3U PD=3U
* device instance $9 r0 *1 9,3.5 NMOS
M$9 10 1 11 11 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $10 r0 *1 12,3.5 NMOS
M$10 11 2 3 11 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS an41

* cell or31$1
* pin VDD
* pin X
* pin C
* pin B
* pin A
* pin VSS
.SUBCKT or31 6 5 4 2 9 3
* net 2 VDD
* net 3 X
* net 4 C
* net 5 B
* net 6 A
* net 9 VSS
* device instance $1 r0 *1 4,23.5 PMOS
M$1 1 6 8 2 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $2 r0 *1 6,23.5 PMOS
M$2 8 5 7 2 PMOS L=1U W=6U AS=3P AD=3P PS=7U PD=7U
* device instance $3 r0 *1 8,23.5 PMOS
M$3 7 4 2 2 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $4 r0 *1 11,23.5 PMOS
M$4 2 1 3 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $5 r0 *1 3,3.5 NMOS
M$5 1 6 9 9 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $6 r0 *1 6,3.5 NMOS
M$6 9 5 1 9 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $7 r0 *1 9,3.5 NMOS
M$7 1 4 9 9 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $8 r0 *1 12,3.5 NMOS
M$8 9 1 3 9 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS or31

* cell nr21$1
* pin X
* pin VDD
* pin A
* pin B
* pin VSS
.SUBCKT nr21 3 4 2 6 1
* net 1 X
* net 2 VDD
* net 3 A
* net 4 B
* net 6 VSS
* device instance $1 r0 *1 3.5,23.5 PMOS
M$1 2 3 5 2 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $2 r0 *1 5.5,23.5 PMOS
M$2 5 4 1 2 PMOS L=1U W=6U AS=3P AD=12P PS=7U PD=16U
* device instance $3 r0 *1 3,3.5 NMOS
M$3 6 3 1 6 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $4 r0 *1 6,3.5 NMOS
M$4 1 4 6 6 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS nr21

* cell na21
* pin X
* pin VDD
* pin B
* pin A
* pin VSS
.SUBCKT na21 4 3 2 6 1
* net 1 X
* net 2 VDD
* net 3 B
* net 4 A
* net 6 VSS
* device instance $1 r0 *1 3,23.5 PMOS
M$1 2 4 1 2 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 6,23.5 PMOS
M$2 1 3 2 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $3 r0 *1 3,3.5 NMOS
M$3 6 4 5 6 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $4 r0 *1 5,3.5 NMOS
M$4 5 3 1 6 NMOS L=1U W=2U AS=1P AD=4P PS=3U PD=8U
.ENDS na21

* cell exor$1
* pin X
* pin VDD
* pin A
* pin B
* pin VSS
.SUBCKT exor 3 4 2 9 1
* net 1 X
* net 2 VDD
* net 3 A
* net 4 B
* net 9 VSS
* device instance $1 r0 *1 11.5,23.5 PMOS
M$1 6 4 2 2 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 14.5,23.5 PMOS
M$2 2 3 6 2 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $3 r0 *1 17.5,23.5 PMOS
M$3 6 5 1 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $4 r0 *1 3,23.5 PMOS
M$4 5 4 7 2 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $5 r0 *1 5,23.5 PMOS
M$5 7 3 2 2 PMOS L=1U W=6U AS=3P AD=12P PS=7U PD=16U
* device instance $6 r0 *1 3,3.5 NMOS
M$6 9 4 5 9 NMOS L=1U W=2U AS=4P AD=2.5P PS=8U PD=4.5U
* device instance $7 r0 *1 6.5,3.5 NMOS
M$7 5 3 9 9 NMOS L=1U W=2U AS=2.5P AD=4P PS=4.5U PD=6U
* device instance $8 r0 *1 11.5,3.5 NMOS
M$8 9 4 8 9 NMOS L=1U W=2U AS=4P AD=1P PS=6U PD=3U
* device instance $9 r0 *1 13.5,3.5 NMOS
M$9 8 3 1 9 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $10 r0 *1 16.5,3.5 NMOS
M$10 1 5 9 9 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS exor

* cell buf8$1
* pin Y
* pin VDD
* pin A
* pin VSS
.SUBCKT buf8 4 3 5 2
* net 2 Y
* net 3 VDD
* net 4 A
* net 5 VSS
* device instance $1 r0 *1 3,23.5 PMOS
M$1 1 4 3 3 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 6,23.5 PMOS
M$2 3 1 2 3 PMOS L=1U W=48U AS=48P AD=54P PS=64U PD=72U
* device instance $10 r0 *1 3,3.5 NMOS
M$10 1 4 5 5 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $11 r0 *1 6,3.5 NMOS
M$11 5 1 2 5 NMOS L=1U W=16U AS=16P AD=18P PS=32U PD=36U
.ENDS buf8

* cell an31$1
* pin Y
* pin VDD
* pin B
* pin A
* pin C
* pin VSS
.SUBCKT an31 5 4 6 2 9 1
* net 1 Y
* net 2 VDD
* net 4 B
* net 5 A
* net 6 C
* net 9 VSS
* device instance $1 r0 *1 3,23.5 PMOS
M$1 3 5 2 2 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 6,23.5 PMOS
M$2 2 4 3 2 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $3 r0 *1 9,23.5 PMOS
M$3 3 6 2 2 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $4 r0 *1 12,23.5 PMOS
M$4 2 3 1 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $5 r0 *1 3,3.5 NMOS
M$5 3 5 8 9 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $6 r0 *1 5,3.5 NMOS
M$6 8 4 7 9 NMOS L=1U W=2U AS=1P AD=1P PS=3U PD=3U
* device instance $7 r0 *1 7,3.5 NMOS
M$7 7 6 9 9 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $8 r0 *1 10,3.5 NMOS
M$8 9 3 1 9 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS an31

* cell sff1m2$1
* pin CK
* pin D
* pin QB
* pin Q
* pin VDD
* pin VSS
.SUBCKT sff1m2 2 4 11 10 9 18 23
* net 2 CK
* net 4 D
* net 9 S
* net 10 QB
* net 11 Q
* net 18 VDD
* net 23 VSS
* device instance $1 r0 *1 12.5,23.5 PMOS
M$1 18 4 19 18 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $2 r0 *1 14.5,23.5 PMOS
M$2 19 1 5 18 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $3 r0 *1 17.5,23.5 PMOS
M$3 5 3 20 18 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $4 r0 *1 19.5,23.5 PMOS
M$4 20 6 18 18 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $5 r0 *1 22.5,23.5 PMOS
M$5 18 5 6 18 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $6 r0 *1 25.5,23.5 PMOS
M$6 6 9 18 18 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $7 r0 *1 28.5,23.5 PMOS
M$7 18 6 21 18 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $8 r0 *1 30.5,23.5 PMOS
M$8 21 3 8 18 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $9 r0 *1 33.5,23.5 PMOS
M$9 8 1 22 18 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $10 r0 *1 35.5,23.5 PMOS
M$10 22 7 18 18 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $11 r0 *1 38.5,23.5 PMOS
M$11 18 8 7 18 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $12 r0 *1 41.5,23.5 PMOS
M$12 7 9 18 18 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $13 r0 *1 49.5,23.5 PMOS
M$13 10 7 18 18 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $14 r0 *1 52.5,23.5 PMOS
M$14 18 10 11 18 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $15 r0 *1 3,23.5 PMOS
M$15 1 2 18 18 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $16 r0 *1 6,23.5 PMOS
M$16 18 1 3 18 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $17 r0 *1 49.5,3.5 NMOS
M$17 10 7 23 23 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $18 r0 *1 52.5,3.5 NMOS
M$18 23 10 11 23 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $19 r0 *1 31,3.5 NMOS
M$19 23 6 15 23 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $20 r0 *1 33,3.5 NMOS
M$20 15 1 8 23 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $21 r0 *1 36,3.5 NMOS
M$21 8 3 16 23 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $22 r0 *1 38,3.5 NMOS
M$22 16 7 23 23 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $23 r0 *1 41,3.5 NMOS
M$23 23 8 17 23 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $24 r0 *1 43,3.5 NMOS
M$24 17 9 7 23 NMOS L=1U W=2U AS=1P AD=4P PS=3U PD=8U
* device instance $25 r0 *1 12.5,3.5 NMOS
M$25 23 4 12 23 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $26 r0 *1 14.5,3.5 NMOS
M$26 12 3 5 23 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $27 r0 *1 17.5,3.5 NMOS
M$27 5 1 13 23 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $28 r0 *1 19.5,3.5 NMOS
M$28 13 6 23 23 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $29 r0 *1 22.5,3.5 NMOS
M$29 23 5 14 23 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $30 r0 *1 24.5,3.5 NMOS
M$30 14 9 6 23 NMOS L=1U W=2U AS=1P AD=4P PS=3U PD=8U
* device instance $31 r0 *1 3,3.5 NMOS
M$31 1 2 23 23 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $32 r0 *1 6,3.5 NMOS
M$32 23 1 3 23 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS sff1m2

* cell or21$1
* pin X
* pin VDD
* pin A
* pin B
* pin VSS
.SUBCKT or21 4 5 2 7 1
* net 1 X
* net 2 VDD
* net 4 A
* net 5 B
* net 7 VSS
* device instance $1 r0 *1 3.5,23.5 PMOS
M$1 3 4 6 2 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $2 r0 *1 5.5,23.5 PMOS
M$2 6 5 2 2 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $3 r0 *1 8.5,23.5 PMOS
M$3 2 3 1 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $4 r0 *1 3,3.5 NMOS
M$4 7 4 3 7 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $5 r0 *1 6,3.5 NMOS
M$5 3 5 7 7 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $6 r0 *1 9,3.5 NMOS
M$6 7 3 1 7 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS or21

* cell na41$1
* pin D
* pin VDD
* pin X
* pin B
* pin A
* pin C
* pin VSS
.SUBCKT na41 5 4 6 1 2 10 3
* net 1 D
* net 2 VDD
* net 3 X
* net 4 B
* net 5 A
* net 6 C
* net 10 VSS
* device instance $1 r0 *1 3,23.5 PMOS
M$1 2 5 3 2 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 6,23.5 PMOS
M$2 3 4 2 2 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $3 r0 *1 9,23.5 PMOS
M$3 2 6 3 2 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $4 r0 *1 12,23.5 PMOS
M$4 3 1 2 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $5 r0 *1 3,3.5 NMOS
M$5 10 5 8 10 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $6 r0 *1 5,3.5 NMOS
M$6 8 4 7 10 NMOS L=1U W=2U AS=1P AD=1P PS=3U PD=3U
* device instance $7 r0 *1 7,3.5 NMOS
M$7 7 6 9 10 NMOS L=1U W=2U AS=1P AD=1P PS=3U PD=3U
* device instance $8 r0 *1 9,3.5 NMOS
M$8 9 1 3 10 NMOS L=1U W=2U AS=1P AD=4P PS=3U PD=8U
.ENDS na41

* cell inv8$1
* pin A
* pin VDD
* pin X
* pin VSS
.SUBCKT inv8 1 2 4 3
* net 1 A
* net 2 VDD
* net 3 X
* net 4 VSS
* device instance $1 r0 *1 3,23.5 PMOS
M$1 2 1 3 2 PMOS L=1U W=48U AS=54P AD=54P PS=72U PD=72U
* device instance $9 r0 *1 3,3.5 NMOS
M$9 4 1 3 4 NMOS L=1U W=16U AS=18P AD=18P PS=36U PD=36U
.ENDS inv8

* cell exnr$1
* pin VDD
* pin X
* pin A
* pin B
* pin VSS
.SUBCKT exnr 3 5 1 9 2
* net 1 VDD
* net 2 X
* net 3 A
* net 5 B
* net 9 VSS
* device instance $1 r0 *1 12.5,23.5 PMOS
M$1 1 5 7 1 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $2 r0 *1 14.5,23.5 PMOS
M$2 7 3 2 1 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $3 r0 *1 17.5,23.5 PMOS
M$3 2 4 1 1 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $4 r0 *1 3,23.5 PMOS
M$4 1 5 4 1 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $5 r0 *1 6,23.5 PMOS
M$5 4 3 1 1 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $6 r0 *1 11.5,3.5 NMOS
M$6 6 5 9 9 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $7 r0 *1 14.5,3.5 NMOS
M$7 9 3 6 9 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $8 r0 *1 17.5,3.5 NMOS
M$8 6 4 2 9 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $9 r0 *1 3,3.5 NMOS
M$9 4 5 8 9 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $10 r0 *1 5,3.5 NMOS
M$10 8 3 9 9 NMOS L=1U W=2U AS=1P AD=4P PS=3U PD=8U
.ENDS exnr

* cell buf4$1
* pin Y
* pin VDD
* pin A
* pin VSS
.SUBCKT buf4 4 3 5 2
* net 2 Y
* net 3 VDD
* net 4 A
* net 5 VSS
* device instance $1 r0 *1 3,23.5 PMOS
M$1 1 4 3 3 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 6,23.5 PMOS
M$2 3 1 2 3 PMOS L=1U W=24U AS=24P AD=30P PS=32U PD=40U
* device instance $6 r0 *1 3,3.5 NMOS
M$6 1 4 5 5 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $7 r0 *1 6,3.5 NMOS
M$7 5 1 2 5 NMOS L=1U W=8U AS=8P AD=10P PS=16U PD=20U
.ENDS buf4

* cell an21$1
* pin VDD
* pin Y
* pin A
* pin B
* pin VSS
.SUBCKT an21 4 5 1 7 3
* net 1 VDD
* net 3 Y
* net 4 A
* net 5 B
* net 7 VSS
* device instance $1 r0 *1 3,23.5 PMOS
M$1 1 4 2 1 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 6,23.5 PMOS
M$2 2 5 1 1 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $3 r0 *1 9,23.5 PMOS
M$3 1 2 3 1 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $4 r0 *1 3,3.5 NMOS
M$4 2 4 6 7 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $5 r0 *1 5,3.5 NMOS
M$5 6 5 7 7 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $6 r0 *1 8,3.5 NMOS
M$6 7 2 3 7 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS an21$1


* cell rff1_r
* pin CK
* pin D
* pin R
* pin QB
* pin Q
* pin VSS
.SUBCKT rff1_r 1 6 13 12 9 2 24
* net 1 CK
* net 2 VDD
* net 6 D
* net 9 R
* net 12 QB
* net 13 Q
* net 24 VSS
* device instance $1 r0 *1 56,23.5 PMOS
M$1 12 10 2 2 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 59,23.5 PMOS
M$2 2 12 13 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $3 r0 *1 37.5,23.5 PMOS
M$3 2 8 21 2 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $4 r0 *1 39.5,23.5 PMOS
M$4 21 5 11 2 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $5 r0 *1 42.5,23.5 PMOS
M$5 11 3 22 2 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $6 r0 *1 44.5,23.5 PMOS
M$6 22 10 2 2 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $7 r0 *1 47.5,23.5 PMOS
M$7 2 11 23 2 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $8 r0 *1 49.5,23.5 PMOS
M$8 23 9 10 2 PMOS L=1U W=6U AS=3P AD=12P PS=7U PD=16U
* device instance $9 r0 *1 19,23.5 PMOS
M$9 2 6 18 2 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $10 r0 *1 21,23.5 PMOS
M$10 18 3 7 2 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $11 r0 *1 24,23.5 PMOS
M$11 7 5 19 2 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $12 r0 *1 26,23.5 PMOS
M$12 19 8 2 2 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $13 r0 *1 29,23.5 PMOS
M$13 2 7 20 2 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $14 r0 *1 31,23.5 PMOS
M$14 20 9 8 2 PMOS L=1U W=6U AS=3P AD=12P PS=7U PD=16U
* device instance $15 r0 *1 9.5,23.5 PMOS
M$15 3 4 2 2 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $16 r0 *1 12.5,23.5 PMOS
M$16 2 3 5 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $17 r0 *1 3,23.5 PMOS
M$17 2 1 4 2 PMOS L=1U W=6U AS=12P AD=12P PS=16U PD=16U
* device instance $18 r0 *1 56,3.5 NMOS
M$18 12 10 24 24 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $19 r0 *1 59,3.5 NMOS
M$19 24 12 13 24 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $20 r0 *1 19,3.5 NMOS
M$20 24 6 14 24 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $21 r0 *1 21,3.5 NMOS
M$21 14 5 7 24 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $22 r0 *1 24,3.5 NMOS
M$22 7 3 15 24 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $23 r0 *1 26,3.5 NMOS
M$23 15 8 24 24 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $24 r0 *1 29,3.5 NMOS
M$24 24 7 8 24 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $25 r0 *1 32,3.5 NMOS
M$25 8 9 24 24 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $26 r0 *1 35,3.5 NMOS
M$26 24 8 16 24 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $27 r0 *1 37,3.5 NMOS
M$27 16 3 11 24 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $28 r0 *1 40,3.5 NMOS
M$28 11 5 17 24 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $29 r0 *1 42,3.5 NMOS
M$29 17 10 24 24 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $30 r0 *1 45,3.5 NMOS
M$30 24 11 10 24 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $31 r0 *1 48,3.5 NMOS
M$31 10 9 24 24 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $32 r0 *1 9.5,3.5 NMOS
M$32 3 4 24 24 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $33 r0 *1 12.5,3.5 NMOS
M$33 24 3 5 24 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $34 r0 *1 3,3.5 NMOS
M$34 24 1 4 24 NMOS L=1U W=2U AS=4P AD=4P PS=8U PD=8U
.ENDS rff1_r

* cell dff1m2_r
* pin CK
* pin D
* pin QB
* pin Q
* pin VSS
.SUBCKT dff1m2_r 1 6 10 9 2 21
* net 1 CK
* net 2 VDD
* net 6 D
* net 9 QB
* net 10 Q
* net 21 VSS
* device instance $1 r0 *1 52,23.5 PMOS
M$1 9 8 2 2 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 55,23.5 PMOS
M$2 2 9 10 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $3 r0 *1 35.5,23.5 PMOS
M$3 2 13 19 2 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $4 r0 *1 37.5,23.5 PMOS
M$4 19 5 14 2 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $5 r0 *1 40.5,23.5 PMOS
M$5 14 3 20 2 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $6 r0 *1 42.5,23.5 PMOS
M$6 20 8 2 2 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $7 r0 *1 45.5,23.5 PMOS
M$7 2 14 8 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $8 r0 *1 19,23.5 PMOS
M$8 2 6 17 2 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $9 r0 *1 21,23.5 PMOS
M$9 17 3 7 2 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $10 r0 *1 24,23.5 PMOS
M$10 7 5 18 2 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $11 r0 *1 26,23.5 PMOS
M$11 18 13 2 2 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $12 r0 *1 29,23.5 PMOS
M$12 2 7 13 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $13 r0 *1 9.5,23.5 PMOS
M$13 3 4 2 2 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $14 r0 *1 12.5,23.5 PMOS
M$14 2 3 5 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $15 r0 *1 3,23.5 PMOS
M$15 2 1 4 2 PMOS L=1U W=6U AS=12P AD=12P PS=16U PD=16U
* device instance $16 r0 *1 52,3.5 NMOS
M$16 9 8 21 21 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $17 r0 *1 55,3.5 NMOS
M$17 21 9 10 21 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $18 r0 *1 35.5,3.5 NMOS
M$18 21 13 16 21 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $19 r0 *1 37.5,3.5 NMOS
M$19 16 3 14 21 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $20 r0 *1 40.5,3.5 NMOS
M$20 14 5 15 21 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $21 r0 *1 42.5,3.5 NMOS
M$21 15 8 21 21 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $22 r0 *1 45.5,3.5 NMOS
M$22 21 14 8 21 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $23 r0 *1 19,3.5 NMOS
M$23 21 6 11 21 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $24 r0 *1 21,3.5 NMOS
M$24 11 5 7 21 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $25 r0 *1 24,3.5 NMOS
M$25 7 3 12 21 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $26 r0 *1 26,3.5 NMOS
M$26 12 13 21 21 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $27 r0 *1 29,3.5 NMOS
M$27 21 7 13 21 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $28 r0 *1 9.5,3.5 NMOS
M$28 3 4 21 21 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $29 r0 *1 12.5,3.5 NMOS
M$29 21 3 5 21 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $30 r0 *1 3,3.5 NMOS
M$30 21 1 4 21 NMOS L=1U W=2U AS=4P AD=4P PS=8U PD=8U
.ENDS dff1m2_r

* cell dff1_r
* pin A,CK
* pin D
* pin QB
* pin Q
* pin VSS
.SUBCKT dff1_r 1 6 11 10 2 21
* net 1 A,CK
* net 2 VDD
* net 6 D
* net 10 QB
* net 11 Q
* net 21 VSS
* device instance $1 r0 *1 52,23.5 PMOS
M$1 10 9 2 2 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 55,23.5 PMOS
M$2 2 10 11 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $3 r0 *1 35.5,23.5 PMOS
M$3 2 8 19 2 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $4 r0 *1 37.5,23.5 PMOS
M$4 19 5 15 2 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $5 r0 *1 40.5,23.5 PMOS
M$5 15 3 20 2 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $6 r0 *1 42.5,23.5 PMOS
M$6 20 9 2 2 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $7 r0 *1 45.5,23.5 PMOS
M$7 2 15 9 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $8 r0 *1 19,23.5 PMOS
M$8 2 6 17 2 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $9 r0 *1 21,23.5 PMOS
M$9 17 3 7 2 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $10 r0 *1 24,23.5 PMOS
M$10 7 5 18 2 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $11 r0 *1 26,23.5 PMOS
M$11 18 8 2 2 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $12 r0 *1 29,23.5 PMOS
M$12 2 7 8 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $13 r0 *1 9.5,23.5 PMOS
M$13 3 4 2 2 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $14 r0 *1 12.5,23.5 PMOS
M$14 2 3 5 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $15 r0 *1 3,23.5 PMOS
M$15 2 1 4 2 PMOS L=1U W=6U AS=12P AD=12P PS=16U PD=16U
* device instance $16 r0 *1 52,3.5 NMOS
M$16 10 9 21 21 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $17 r0 *1 55,3.5 NMOS
M$17 21 10 11 21 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $18 r0 *1 35.5,3.5 NMOS
M$18 21 8 14 21 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $19 r0 *1 37.5,3.5 NMOS
M$19 14 3 15 21 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $20 r0 *1 40.5,3.5 NMOS
M$20 15 5 16 21 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $21 r0 *1 42.5,3.5 NMOS
M$21 16 9 21 21 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $22 r0 *1 45.5,3.5 NMOS
M$22 21 15 9 21 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $23 r0 *1 19,3.5 NMOS
M$23 21 6 12 21 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $24 r0 *1 21,3.5 NMOS
M$24 12 5 7 21 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $25 r0 *1 24,3.5 NMOS
M$25 7 3 13 21 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $26 r0 *1 26,3.5 NMOS
M$26 13 8 21 21 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $27 r0 *1 29,3.5 NMOS
M$27 21 7 8 21 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $28 r0 *1 9.5,3.5 NMOS
M$28 3 4 21 21 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $29 r0 *1 12.5,3.5 NMOS
M$29 21 3 5 21 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $30 r0 *1 3,3.5 NMOS
M$30 21 1 4 21 NMOS L=1U W=2U AS=4P AD=4P PS=8U PD=8U
.ENDS dff1_r

* cell sff1m2_r
* pin CK
* pin D
* pin S
* pin QB
* pin Q
* pin VSS
.SUBCKT sff1m2_r 1 5 12 11 10 19 24
* net 1 CK
* net 5 D
* net 10 S
* net 11 QB
* net 12 Q
* net 19 VDD
* net 24 VSS
* device instance $1 r0 *1 56,23.5 PMOS
M$1 11 8 19 19 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 59,23.5 PMOS
M$2 19 11 12 19 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $3 r0 *1 19,23.5 PMOS
M$3 19 5 20 19 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $4 r0 *1 21,23.5 PMOS
M$4 20 2 6 19 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $5 r0 *1 24,23.5 PMOS
M$5 6 4 21 19 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $6 r0 *1 26,23.5 PMOS
M$6 21 7 19 19 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $7 r0 *1 29,23.5 PMOS
M$7 19 6 7 19 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $8 r0 *1 32,23.5 PMOS
M$8 7 10 19 19 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $9 r0 *1 35,23.5 PMOS
M$9 19 7 22 19 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $10 r0 *1 37,23.5 PMOS
M$10 22 4 9 19 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $11 r0 *1 40,23.5 PMOS
M$11 9 2 23 19 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $12 r0 *1 42,23.5 PMOS
M$12 23 8 19 19 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $13 r0 *1 45,23.5 PMOS
M$13 19 9 8 19 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $14 r0 *1 48,23.5 PMOS
M$14 8 10 19 19 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $15 r0 *1 9.5,23.5 PMOS
M$15 2 3 19 19 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $16 r0 *1 12.5,23.5 PMOS
M$16 19 2 4 19 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $17 r0 *1 3,23.5 PMOS
M$17 19 1 3 19 PMOS L=1U W=6U AS=12P AD=12P PS=16U PD=16U
* device instance $18 r0 *1 56,3.5 NMOS
M$18 11 8 24 24 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $19 r0 *1 59,3.5 NMOS
M$19 24 11 12 24 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $20 r0 *1 37.5,3.5 NMOS
M$20 24 7 16 24 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $21 r0 *1 39.5,3.5 NMOS
M$21 16 2 9 24 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $22 r0 *1 42.5,3.5 NMOS
M$22 9 4 17 24 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $23 r0 *1 44.5,3.5 NMOS
M$23 17 8 24 24 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $24 r0 *1 47.5,3.5 NMOS
M$24 24 9 18 24 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $25 r0 *1 49.5,3.5 NMOS
M$25 18 10 8 24 NMOS L=1U W=2U AS=1P AD=4P PS=3U PD=8U
* device instance $26 r0 *1 19,3.5 NMOS
M$26 24 5 13 24 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $27 r0 *1 21,3.5 NMOS
M$27 13 4 6 24 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $28 r0 *1 24,3.5 NMOS
M$28 6 2 15 24 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $29 r0 *1 26,3.5 NMOS
M$29 15 7 24 24 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $30 r0 *1 29,3.5 NMOS
M$30 24 6 14 24 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $31 r0 *1 31,3.5 NMOS
M$31 14 10 7 24 NMOS L=1U W=2U AS=1P AD=4P PS=3U PD=8U
* device instance $32 r0 *1 9.5,3.5 NMOS
M$32 2 3 24 24 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $33 r0 *1 12.5,3.5 NMOS
M$33 24 2 4 24 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $34 r0 *1 3,3.5 NMOS
M$34 24 1 3 24 NMOS L=1U W=2U AS=4P AD=4P PS=8U PD=8U
.ENDS sff1m2_r

* cell sff1_r
* pin CK
* pin D
* pin S
* pin QB
* pin Q
* pin VSS
.SUBCKT sff1_r 1 6 13 12 11 2 24
* net 1 CK
* net 2 VDD
* net 6 D
* net 11 S
* net 12 QB
* net 13 Q
* net 24 VSS
* device instance $1 r0 *1 56,23.5 PMOS
M$1 12 10 2 2 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 59,23.5 PMOS
M$2 2 12 13 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $3 r0 *1 19,23.5 PMOS
M$3 2 6 20 2 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $4 r0 *1 21,23.5 PMOS
M$4 20 3 7 2 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $5 r0 *1 24,23.5 PMOS
M$5 7 5 21 2 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $6 r0 *1 26,23.5 PMOS
M$6 21 8 2 2 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $7 r0 *1 29,23.5 PMOS
M$7 2 7 8 2 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $8 r0 *1 32,23.5 PMOS
M$8 8 11 2 2 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $9 r0 *1 35,23.5 PMOS
M$9 2 8 22 2 PMOS L=1U W=6U AS=6P AD=7.5P PS=8U PD=8.5U
* device instance $10 r0 *1 38.5,23.5 PMOS
M$10 22 5 9 2 PMOS L=1U W=6U AS=7.5P AD=6P PS=8.5U PD=8U
* device instance $11 r0 *1 41.5,23.5 PMOS
M$11 9 3 23 2 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $12 r0 *1 43.5,23.5 PMOS
M$12 23 10 2 2 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $13 r0 *1 46.5,23.5 PMOS
M$13 2 9 10 2 PMOS L=1U W=6U AS=6P AD=6P PS=8U PD=8U
* device instance $14 r0 *1 49.5,23.5 PMOS
M$14 10 11 2 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $15 r0 *1 9.5,23.5 PMOS
M$15 3 4 2 2 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $16 r0 *1 12.5,23.5 PMOS
M$16 2 3 5 2 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $17 r0 *1 3,23.5 PMOS
M$17 2 1 4 2 PMOS L=1U W=6U AS=12P AD=12P PS=16U PD=16U
* device instance $18 r0 *1 56,3.5 NMOS
M$18 12 10 24 24 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $19 r0 *1 59,3.5 NMOS
M$19 24 12 13 24 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $20 r0 *1 37.5,3.5 NMOS
M$20 24 8 18 24 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $21 r0 *1 39.5,3.5 NMOS
M$21 18 3 9 24 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $22 r0 *1 42.5,3.5 NMOS
M$22 9 5 17 24 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $23 r0 *1 44.5,3.5 NMOS
M$23 17 10 24 24 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $24 r0 *1 47.5,3.5 NMOS
M$24 24 9 19 24 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $25 r0 *1 49.5,3.5 NMOS
M$25 19 11 10 24 NMOS L=1U W=2U AS=1P AD=4P PS=3U PD=8U
* device instance $26 r0 *1 19,3.5 NMOS
M$26 24 6 14 24 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $27 r0 *1 21,3.5 NMOS
M$27 14 5 7 24 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $28 r0 *1 24,3.5 NMOS
M$28 7 3 15 24 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $29 r0 *1 26,3.5 NMOS
M$29 15 8 24 24 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $30 r0 *1 29,3.5 NMOS
M$30 24 7 16 24 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $31 r0 *1 31,3.5 NMOS
M$31 16 11 8 24 NMOS L=1U W=2U AS=1P AD=4P PS=3U PD=8U
* device instance $32 r0 *1 9.5,3.5 NMOS
M$32 3 4 24 24 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $33 r0 *1 12.5,3.5 NMOS
M$33 24 3 5 24 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $34 r0 *1 3,3.5 NMOS
M$34 24 1 4 24 NMOS L=1U W=2U AS=4P AD=4P PS=8U PD=8U
.ENDS sff1_r

* cell rff1m2_r
* pin Q
* pin CK
* pin D
* pin R
* pin QB
* pin VSS
.SUBCKT rff1m2_r 2 7 1 12 10 3 24
* net 1 Q
* net 2 CK
* net 3 VDD
* net 7 D
* net 10 R
* net 12 QB
* net 24 VSS
* device instance $1 r0 *1 56,23.5 PMOS
M$1 12 11 3 3 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 59,23.5 PMOS
M$2 3 12 1 3 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $3 r0 *1 37.5,23.5 PMOS
M$3 3 9 21 3 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $4 r0 *1 39.5,23.5 PMOS
M$4 21 6 15 3 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $5 r0 *1 42.5,23.5 PMOS
M$5 15 4 22 3 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $6 r0 *1 44.5,23.5 PMOS
M$6 22 11 3 3 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $7 r0 *1 47.5,23.5 PMOS
M$7 3 15 23 3 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $8 r0 *1 49.5,23.5 PMOS
M$8 23 10 11 3 PMOS L=1U W=6U AS=3P AD=12P PS=7U PD=16U
* device instance $9 r0 *1 19,23.5 PMOS
M$9 3 7 18 3 PMOS L=1U W=6U AS=12P AD=3P PS=16U PD=7U
* device instance $10 r0 *1 21,23.5 PMOS
M$10 18 4 8 3 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $11 r0 *1 24,23.5 PMOS
M$11 8 6 19 3 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $12 r0 *1 26,23.5 PMOS
M$12 19 9 3 3 PMOS L=1U W=6U AS=3P AD=6P PS=7U PD=8U
* device instance $13 r0 *1 29,23.5 PMOS
M$13 3 8 20 3 PMOS L=1U W=6U AS=6P AD=3P PS=8U PD=7U
* device instance $14 r0 *1 31,23.5 PMOS
M$14 20 10 9 3 PMOS L=1U W=6U AS=3P AD=12P PS=7U PD=16U
* device instance $15 r0 *1 9.5,23.5 PMOS
M$15 4 5 3 3 PMOS L=1U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $16 r0 *1 12.5,23.5 PMOS
M$16 3 4 6 3 PMOS L=1U W=6U AS=6P AD=12P PS=8U PD=16U
* device instance $17 r0 *1 3,23.5 PMOS
M$17 3 2 5 3 PMOS L=1U W=6U AS=12P AD=12P PS=16U PD=16U
* device instance $18 r0 *1 56,3.5 NMOS
M$18 12 11 24 24 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $19 r0 *1 59,3.5 NMOS
M$19 24 12 1 24 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $20 r0 *1 19,3.5 NMOS
M$20 24 7 13 24 NMOS L=1U W=2U AS=4P AD=1P PS=8U PD=3U
* device instance $21 r0 *1 21,3.5 NMOS
M$21 13 6 8 24 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $22 r0 *1 24,3.5 NMOS
M$22 8 4 14 24 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $23 r0 *1 26,3.5 NMOS
M$23 14 9 24 24 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $24 r0 *1 29,3.5 NMOS
M$24 24 8 9 24 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $25 r0 *1 32,3.5 NMOS
M$25 9 10 24 24 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $26 r0 *1 35,3.5 NMOS
M$26 24 9 16 24 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $27 r0 *1 37,3.5 NMOS
M$27 16 4 15 24 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $28 r0 *1 40,3.5 NMOS
M$28 15 6 17 24 NMOS L=1U W=2U AS=2P AD=1P PS=4U PD=3U
* device instance $29 r0 *1 42,3.5 NMOS
M$29 17 11 24 24 NMOS L=1U W=2U AS=1P AD=2P PS=3U PD=4U
* device instance $30 r0 *1 45,3.5 NMOS
M$30 24 15 11 24 NMOS L=1U W=2U AS=2P AD=2P PS=4U PD=4U
* device instance $31 r0 *1 48,3.5 NMOS
M$31 11 10 24 24 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $32 r0 *1 9.5,3.5 NMOS
M$32 4 5 24 24 NMOS L=1U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $33 r0 *1 12.5,3.5 NMOS
M$33 24 4 6 24 NMOS L=1U W=2U AS=2P AD=4P PS=4U PD=8U
* device instance $34 r0 *1 3,3.5 NMOS
M$34 24 2 5 24 NMOS L=1U W=2U AS=4P AD=4P PS=8U PD=8U
.ENDS rff1m2_r


